library IEEE; use IEEE.STD_LOGIC_1164.all;
entity rom is
port
(
adr: in STD_LOGIC_VECTOR(1 downto 0);
dout: out STD_LOGIC_VECTOR(2 downto 0)
);
end;
architecture synth of rom is
begin
--process(all) begin--VHDL2008
process (adr) begin
case adr is
when "00" => dout <= "011";
when "01" => dout <= "110";
when "10" => dout <= "100";
when "11" => dout <= "010";
end case;
end process;
end;
